module MUL_datapath(eqz, LdA, LdB, LdP, clrP, decB, data_in, clk);

	input LdA, LdB, LdP, clrP, decB, clk;
	input [15:0] data_in;
	output eqz;
	wire [15:0] X, Y, Z, Bout, Bus;

	PIPO1 A(X, Bus, LdA, clk);
	PIPO2 P(Y, Z, LdP, clrP, clk);
	CNTR B(Bout, Bus, LdB, decB, clk);
	ADD AD(Z, X, Y);
	EQZ COMP(eqz, Bout);

endmodule

module PIPO1(dout, din, ld, clk);

	input [15:0] din;
	input ld, clk;
	output reg[15:0] dout;

	always @(posedge clk)
		if(ld) dout <= din;

endmodule

module PIPO2(dout, in, ld, clr, clk);

	input [15:0] din;
	input ld, clr, clk;
	output reg [15:0] dout;

	always @(posedge clk) begin
		if(clr) dout <= 16'b0;
		else if (ld) dout <= din;
	end

endmodule
